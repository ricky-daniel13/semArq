`timescale 1ns/1ns
module actividad03_tb();
reg entrada1; reg entrada2; output salidaand;
wire salidaand; wire salidaor; wire salidaxor; wire salidanot; wire salidanand; wire salidayes; wire salidanor; wire salidaxnor );
actividad03 a(
reg.(reg),
entrada1.(entrada1),
reg.(reg),
entrada2.(entrada2),
output.(output),
salidaand.(salidaand),
wire.(wire),
salidaand.(salidaand),
wire.(wire),
salidaor.(salidaor),
wire.(wire),
salidaxor.(salidaxor),
wire.(wire),
salidanot.(salidanot),
wire.(wire),
salidanand.(salidanand),
wire.(wire),
salidayes.(salidayes),
wire.(wire),
salidanor.(salidanor),
wire.(wire),
salidaxnor.(salidaxnor),
).()),
);
initial
begin
end
endmodule
