module rom(
	input [4:0]dir,
	output reg [31:0]inst
);
reg [7:0] isa [0:25];
always @*
begin
	
end
endmodule