module memorias(
	input 
		en,
		clk,
	input [4:0]dir,
	input [7:0]dataIn,
	output reg [7:0]dataOut
);
endmodule